library ieee;
use ieee.std_logic_1164.all;

entity riscy_top is
    port(
        clk : in std_logic;
        reset : in std_logic
    );
end entity;

architecture behav of riscy_top is
begin
end architecture;